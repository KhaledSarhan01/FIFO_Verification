import shared_pkg::*;

module FIFO_tb(FIFO_if.TEST if_handle);
    
endmodule