import shared_pkg::*;

module FIFO_MONITOR(FIFO_if.MONITPR if_handle);
    
endmodule