import shared_pkg::*;

module FIFO_MONITOR(FIFO_if.MONITOR if_handle);
    
endmodule